`timescale 1ns / 1ps

module hex7seg(
    input [3:0] n,
    output [6:0] seg
    );   
   assign seg[0] = (~n[3]&~n[2]&~n[1]&n[0]) |(~n[3]&n[2]&~n[1]&~n[0]) | (n[3]&~n[2]&n[1]&n[0]) |(n[3]&n[2]&~n[1]&n[0]);
   assign seg[1] = (~n[3]&n[2]&~n[1]&n[0]) |(~n[3]&n[2]&n[1]&~n[0]) |(n[3]&~n[2]&n[1]&n[0]) |(n[3]&n[2]&~n[1]&~n[0]) |(n[3]&n[2]&n[1]&~n[0]) |(n[3]&n[2]&n[1]&n[0]);
   assign seg[2] = (~n[3]&~n[2]&n[1]&~n[0]) |(n[3]&n[2]&~n[1]&~n[0]) |(n[3]&n[2]&n[1]&~n[0]) |(n[3]&n[2]&n[1]&n[0]);
   assign seg[3] = (~n[3]&~n[2]&~n[1]&n[0]) |(~n[3]&n[2]&~n[1]&~n[0]) |(~n[3]&n[2]&n[1]&n[0]) |(n[3]&~n[2]&~n[1]&n[0]) |(n[3]&~n[2]&n[1]&~n[0]) |(n[3]&n[2]&n[1]&n[0]);
   assign seg[4] = (~n[3]&~n[2]&~n[1]&n[0]) |(~n[3]&~n[2]&n[1]&n[0]) |(~n[3]&n[2]&~n[1]&~n[0]) |(~n[3]&n[2]&~n[1]&n[0]) |(~n[3]&n[2]&n[1]&n[0]) |(n[3]&~n[2]&~n[1]&n[0]);
   assign seg[5] = (~n[3]&~n[2]&~n[1]&n[0]) |(~n[3]&~n[2]&n[1]&~n[0]) |(~n[3]&~n[2]&n[1]&n[0]) |(~n[3]&n[2]&n[1]&n[0]) |(n[3]&n[2]&~n[1]&n[0]);
   assign seg[6] = (~n[3]&~n[2]&~n[1]&~n[0]) |(~n[3]&~n[2]&~n[1]&n[0]) |(~n[3]&n[2]&n[1]&n[0]) |(n[3]&n[2]&~n[1]&~n[0]);
endmodule
/*
1
(~n[3]&~n[2]&~n[1]&~n[0]) |
2
(~n[3]&~n[2]&~n[1]&n[0]) |
3
(~n[3]&~n[2]&n[1]&~n[0]) |
4
(~n[3]&~n[2]&n[1]&n[0]) |
5
(~n[3]&n[2]&~n[1]&~n[0]) |
6
(~n[3]&n[2]&~n[1]&n[0]) |
7
(~n[3]&n[2]&n[1]&~n[0]) |
8
(~n[3]&n[2]&n[1]&n[0]) |
9
(n[3]&~n[2]&~n[1]&~n[0]) |
10
(n[3]&~n[2]&~n[1]&n[0]) |
11
(n[3]&~n[2]&n[1]&~n[0]) |
12
(n[3]&~n[2]&n[1]&n[0]) |
13
(n[3]&n[2]&~n[1]&~n[0]) |
14
(n[3]&n[2]&~n[1]&n[0]) |
15
(n[3]&n[2]&n[1]&~n[0]) |
16
(n[3]&n[2]&n[1]&n[0]) |
*/

